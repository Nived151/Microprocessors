module data_mem();
input address_bus[0:7];
input data_in[0:7];
reg data_out[0:7];
input r_w;

endmodule