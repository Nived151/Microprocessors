module program_mem();
input program_mem_address_bus[0:7];
output program_mem_data_out[0:16];
reg op_codes[5:0];




endmodule