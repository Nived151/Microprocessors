module program_mem();
input program_mem_address_bus[0:7];
reg program_mem_data_out[0:15];

endmodule